module chessEngine(

);



endmodule
